module NotBinario(in,out);
	input in;
	output out;
	
	NandBinario n(in,in,out);
endmodule
	
